* File: inversorp4.pex.netlist
* Created: Tue Jul  4 17:33:46 2023
* Program "Calibre xRC"
* Version "v2006.2_16.16"
* 
.subckt INVERSORP4 OUT IN VSS VDD
mM0 VSS IN OUT VSS NMOS4 L=3.5e-07 W=4e-06 AD=3.8e-12 AS=3.4e-12 PD=5.9e-06
+ PS=5.7e-06 NRD=0.10625 NRS=0.10625
mM1 VDD IN OUT VDD PMOS4 L=3.5e-07 W=1.175e-05 AD=1.11625e-11 AS=9.9875e-12
+ PD=1.365e-05 PS=1.345e-05 NRD=0.0361702 NRS=0.0361702
*
.include "inversorp4.pex.netlist.INVERSORP4.pxi"
*
.ends
*
*
